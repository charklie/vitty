module ascii_logos

const orange = '\u001b[31;1m'
const lightblue = '\u001b[36;1m'
const blue = '\u001b[34m'
const white = '\u001b[37m'
const reset = '\u001b[0m'

pub const windows11_logo = '
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}

${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}
${blue}################  ################${reset}'

pub const windows10_logo = '
${blue}                                ..,${reset}
${blue}                    ....,,:;+ccllll${reset}
${blue}      ...,,+:;  cllllllllllllllllll${reset}
${blue},cclllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}

${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}llllllllllllll  lllllllllllllllllll${reset}
${blue}`\'ccllllllllll  lllllllllllllllllll${reset}
${blue}       `\' \\*::  :ccllllllllllllllll${reset}
${blue}                       ````\'\'*::cll${reset}
${blue}                                  `${reset}'

pub const ubuntu_logo = '
${orange}            .-/+oossssoo+\\-.${reset}
${orange}       ´:+ssssssssssssssssss+:`${reset}
${orange}     -+ssssssssssssssssssyyssss+-${reset}
${orange}   .ossssssssssssssssss${white}dMMMNy${orange}sssso.${reset}
${orange}   /sssssssssss${white}hdmmNNmmyNMMMMh${orange}ssssss\\${reset}
${orange}  +sssssssss${white}hm${orange}yd${white}MMMMMMMNddddy${orange}ssssssss+${reset}
${orange} /ssssssss${white}hNMMM${orange}yh${white}hyyyyhmNMMMNh${orange}ssssssss\\${reset}
${orange}.ssssssss${white}dMMMNh${orange}ssssssssss${white}hNMMMd${orange}ssssssss.${reset}
${orange}+ssss${white}hhhyNMMNy${orange}ssssssssssss${white}yNMMMy${orange}sssssss+${reset}
${orange}oss${white}yNMMMNyMMh${orange}ssssssssssssss${white}hmmmh${orange}ssssssso${reset}
${orange}oss${white}yNMMMNyMMh${orange}sssssssssssssshmmmh${orange}ssssssso${reset}
${orange}+ssss${white}hhhyNMMNy${orange}ssssssssssss${white}yNMMMy${orange}sssssss+${reset}
${orange}.ssssssss${white}dMMMNh${orange}ssssssssss${white}hNMMMd${orange}ssssssss.${reset}
${orange} \\ssssssss${white}hNMMM${orange}yh${white}hyyyyhdNMMMNh${orange}ssssssss/${reset}
${orange}  +sssssssss${white}dm${orange}yd${white}MMMMMMMMddddy${orange}ssssssss+${reset}
${orange}   \\sssssssssss${white}hdmNNNNmyNMMMMh${orange}ssssss/${reset}
${orange}    .ossssssssssssssssss${white}dMMMNy${orange}sssso.${reset}
${orange}      -+sssssssssssssssss${white}yyy${orange}ssss+-${reset}
${orange}        `:+ssssssssssssssssss+:`${reset}
${orange}            .-\\+oossssoo+/-.${reset}'

pub const arch_logo = '
${lightblue}                   -`${reset}
${lightblue}                  .o+`${reset}
${lightblue}                 `ooo/${reset}
${lightblue}                `+oooo:${reset}
${lightblue}               `+oooooo:${reset}
${lightblue}               -+oooooo+:${reset}
${lightblue}             `/:-:++oooo+:${reset}
${lightblue}            `/++++/+++++++:${reset}
${lightblue}           `/++++++++++++++:${reset}
${lightblue}          `/+++ooooooooooooo/`${reset}
${lightblue}         ./ooosssso++osssssso+`${reset}
${lightblue}        .oossssso-````/ossssss+`${reset}
${lightblue}       -osssssso.      :ssssssso.${reset}
${lightblue}      :osssssss/        osssso+++.${reset}
${lightblue}     /ossssssss/        +ssssooo/-${reset}
${lightblue}   `/ossssso+/:-        -:/+osssso+-${reset}
${lightblue}  `+sso+:-`                 `.-/+oso:${reset}
${lightblue} `++:.                           `-/+/${reset}
${lightblue} .`                                 `/.${reset}'
