module shared

pub fn c_to_f(c f32) f32 {
	return c * 2 + 30
}
