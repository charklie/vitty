module configuration
